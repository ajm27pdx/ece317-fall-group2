i   ����MbP?���ư>                ��         ����MbP?���ư>      �?                          !         �?2                 I1      I1      H   �       	           6                 VP1     I01     �   �      -C��6?2                 C1  �@� C1      �   �           
           6                 IP1     V01     �   �              �                 GND1            H   0      {�G�z�?2                 R1      R1      x  �                      �                 MOD1            �  �         �               @              �?           �                  CLK1              �           �y�Cn�+?           2   	              SW1     S1      x  �                  �   
   H     H   (                            �      H   �   H   �                             �      H   �   �   �                             �      �   �   �   �                             �      �   �   �   �                              �      x     x                              �      �     x                              �      �     �                                �      H     �                                �      �   �   x  �                              �      x  �   x  �                             �      x  �   x  �                             �      (  �   h  �                              �      �  �   �  �                              �      �  �   �                              �      �    �                               �      �  �   �                              �      �   p   �  p                              �      �   p   �   �                     