i   ���Q��?H����׊>                ��         ���Q��?���ư>      �?                             ���מYB?2                  L1 E1   L1  	�  �                     9@2                 R1  @� R1      P  �              -C��6?2                 C1 j@c?jC1 j@c?j   �           	           6                 VP2     I01     �  �   	           6                 VP1     I02     @  �             $@2                 V1  r  V1   F (   �                  2                 SW2 �c�tS1      �   �                  �   	   �   @   �   @                             �      �   �   �   �                             �      X   �   �   �                              2                 SW3     S2      �   @                 �      X   @   �   @                              �                 CLK1            �   �   �����>�h㈵��>           �                  CLK2            H   �           �h㈵��>           �      X   @   X   �                             �      X   �   X   �                             �      �   @   �   �                            �      �   �   �   �                            �      �  �   �  �                             �      P  �   P  �                             �      P  �   �  �                             �   
      �      �                             �         �   P  �                             �      �   �   �   �                             �      @  �   @  �                             �      �   �   @  �                             �      @  �      �                             �      �  �   �  �                             �      P  �   P  �                             �   !   P  �   �  �                             �         �      �                             �   "   �  �      �                             �   #      �   P  �                             �   $   @  �   @  �                             �   %   (   (   (   �                             �   &   (   (   �   (                             �   (   �   �   @  �                             �   )   @  �   �  �                             �       �   X   �   �                            �   *   �   �   �   �                            �   '              GND1  s   e s   `   �              �   +   (   �   `   �                             �   ,   `   �   �   �                     