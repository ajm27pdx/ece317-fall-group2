i   ���Q��?H����׊>                ��         ���Q��?���ư>      �?                             ���מYB?2                  L1 E1   L1  	  �                     9@2                 R1  @� R1      �  �              -C��6?2                 C1 j@c?jC1 j@c?jh  �           	           6                 VP2     I01        �   	           6                 VP1     I02     �  �             $@2                 V1  r  V1   F (   �                  2                 SW2 �c�tS1      �   �                  �   	   �   @   �   @                             �      �   �   �   �                             �      X   �   �   �                              2                 SW3     S2      �   @                 �      X   @   �   @                              �                  CLK2            H   �           -C��6�>           �      X   @   X   �                             �      X   �   X   �                             �      �   �   �   �                            �         �      �                             �      �  �   �  �                             �      �  �      �                             �   
   h  �   h  �                             �      h  �   �  �                             �      �   �   �   �                             �      �  �   �  �                             �      �  �   h  �                             �         �      �                             �      �  �   �  �                             �   !   �  �      �                             �      h  �   h  �                             �   "      �   h  �                             �   #   h  �   �  �                             �   $   �  �   �  �                             �   %   (   (   (   �                             �   &   (   (   �   (                             �   )   �  �   �  �                             �       �   H   �   x                             �   *   �   �   �   �                            �   '              GND1  s   e s   `   �              �   +   (   �   `   �                             �   ,   `   �   �   �                          jA�                 MOD1 �ʂ �L�u�L@  �         �?                      @-C��6�>          @2                 V2 �  V2     �   �                  �      �   x   �   x                              �   (   �   X   �   x                            �   -   �   x   �   �                            �   .   �   H   �  H                              �   0   �   p     p                              �   1   �   p   �   x                             �   /   �  H   �  �                             �   3   h  X   h  �                              �   4   �   X   h  X                              �   5   �   X   �   �                             �   6   �   �   �   �                              �   7   �   @   �   �                            �   8   �   �   �   �                            �      �   �   �   �                             �   9   �   �   �   �                             �   :   �   �   �  �                     